
class empty_executor_trait_s extends executor_trait_s;
endclass
