
typedef class object_c;
typedef class object_ref_c;

class input_c #(type T=object_c) extends object_ref_c #(T);

    function new();
        super.new();
    endfunction


endclass