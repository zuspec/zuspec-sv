
class executor_trait_s extends empty_executor_trait_s;
endclass

