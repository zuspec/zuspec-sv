
typedef component_c component_queue_h[$];
typedef class pool_c;

class component_c extends typed_obj_c;
    int                     comp_id;
    string                  name;
    component_c             parent;
    
    pool_c                pool_m;


    /**
     * Map of component type to list of component instances
     * at this level and below.
     */
    component_queue_h       comp_t_inst_m[obj_type_c];


    // Each component needs a map of action-claim refs to pool
    executor_base  executor_m[];

    // aspace_t_map
    // executor_t_map

    function new(string name, component_ctor_ctxt ctxt, component_c parent=null);
        $display("component_c::new: %0s ctxt=%p", name, ctxt);
        this.name = name;
        this.parent = parent;
        if (ctxt != null) begin
            this.comp_id = ctxt.actor.comp_l.size();
            ctxt.actor.comp_l.push_back(this);
        end else begin
            this.comp_id = -1;
        end
    endfunction

    /**
     * Adds a component instance to the map of comp_t -> [comp_inst] map
     */
    function void add_comp_inst(component_c comp);
        obj_type_c comp_t = comp.get_obj_type();
        $display("add_comp_inst: %0s (%0s)", comp.name, this.name);
        $display("comp_obj_type: %0p", comp_t);
        if (comp_t_inst_m.exists(comp_t)) begin
            comp_t_inst_m[comp_t].push_back(comp);
        end else begin
            component_queue_h l;
            l.push_back(comp);
            comp_t_inst_m[comp_t] = l;
        end
        $display("Contains: %0d", comp_t_inst_m[comp_t].size);
    endfunction

    virtual function void init_down(executor_base exec_b);
    endfunction

    virtual function void init(executor_base exec_b);
    endfunction

    virtual function void init_up(executor_base exec_b);
    endfunction

    virtual function void start(executor_base exec_b);
    endfunction

    virtual function bit check();
        return 1;
    endfunction

    virtual function actor_c get_actor();
        component_c c = parent;
        actor_c actor;

        while (c.parent != null) begin
            c = c.parent;
        end
        $cast(actor, c);
        return actor;
    endfunction

    virtual function executor_base get_default_executor();
        component_c c = parent;
        actor_c actor;

        while (c.parent != null) begin
            c = c.parent;
        end
        $cast(actor, c);
        return actor.get_default_executor();
    endfunction

endclass
