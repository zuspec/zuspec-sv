
class addr_trait_s;
endclass
