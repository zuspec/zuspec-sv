
class transparent_addr_region_s extends addr_region_s;

    static function transparent_addr_region_s create_default();
        transparent_addr_region_s ret = new();
        return ret;
    endfunction

endclass