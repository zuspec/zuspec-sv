typedef class solve_pool_c;

class solve_resource_pool_c extends solve_pool_c;
    bit[31:0]               size;
endclass