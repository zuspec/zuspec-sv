
class empty_executor_trait_s extends object;
endclass
