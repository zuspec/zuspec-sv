
class solve_pool_c;
endclass
