
class flow_obj_pool_c;
endclass

