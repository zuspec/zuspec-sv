
class addr_region_s extends addr_region_base_s;
    bit[31:0]   size;
endclass
