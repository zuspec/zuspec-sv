
class addr_claim_base_s;
endclass
