
typedef class storage_handle_c; 

class addr_claim_base_s extends object_ref_c #(storage_handle_c);
    function new();
        super.new();
    endfunction

endclass
