
typedef class object_refcnt_c;

class object_mgr_c;

    virtual function void release_obj(object_refcnt_c obj);
    endfunction

endclass
