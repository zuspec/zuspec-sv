typedef class activity_ctxt_c;

class activity_builder_c;
    virtual function void build(activity_ctxt_c ctxt);
    endfunction

endclass