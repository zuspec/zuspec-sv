
typedef class pool_c;

class flow_obj_c extends object;
    pool_c      pool;
endclass

