
class obj_type_c;
    string  name;

    function new(string name);
        this.name = name;
    endfunction

    static function obj_type_c get_type();
    endfunction

endclass
