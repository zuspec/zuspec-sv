
class solve_traversal_context_c;
    action_type_c                 action_t;
    rand bit[31:0]                comp_id;
    bit[31:0]                     comp_id_l[$];
    rand pool_ref_c               pool_refs_l[$];
endclass