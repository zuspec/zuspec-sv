
class storage_handle_s extends object_pool_base;
    bit[63:0]           addr;

endclass