
class solve_compset_c;
    bit[31:0]            comp_id_l[$];
endclass