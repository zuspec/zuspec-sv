
typedef class obj_type_c;

class typed_obj_c;

    static function obj_type_c get_type();
        return null;
    endfunction

endclass
