
typedef class object_c;

class executor_trait_s extends object_c;
endclass

