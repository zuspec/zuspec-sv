
class solve_pool2comp_map_c;
    bit[31:0]               pool2comp_m[$];
endclass
