
class executor_trait_s extends object;
endclass

