
class empty_executor_trait_s extends object;
    `zsp_typed_obj_util(empty_executor_trait_s)
endclass
