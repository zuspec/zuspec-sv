
class solve_pool_ref_c;
    rand bit[31:0]          pool_id;
    pool_base_c             pools[$];
endclass
