
class activity_par_c extends activity_c;
    activity_c      sub_activities[$];

    function new(actor_c actor);
        super.new(actor);s
    endfunction


endclass
