
typedef class object_c;

class empty_executor_trait_s extends object_c;
    `zsp_typed_obj_util(empty_executor_trait_s)
endclass
