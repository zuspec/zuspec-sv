/*
 * activity_ctxt_seq_c.svh
 *
 * Copyright 2023 Matthew Ballance and Contributors
 *
 * Licensed under the Apache License, Version 2.0 (the "License"); you may 
 * not use this file except in compliance with the License.  
 * You may obtain a copy of the License at:
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software 
 * distributed under the License is distributed on an "AS IS" BASIS, 
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.  
 * See the License for the specific language governing permissions and 
 * limitations under the License.
 *
 * Created on:
 *     Author:
 */

typedef class activity_ctxt_c;

class activity_ctxt_seq_c extends activity_ctxt_c;

    function new(activity_ctxt_c parent);
        super.new(parent);
    endfunction

    virtual task add(activity_c activity);
        activity.run(this);
    endtask

    static function activity_ctxt_seq_c mk(activity_ctxt_c parent);
        activity_ctxt_seq_c ctxt = new(parent);
        return ctxt;
    endfunction

endclass

