typedef class object;
typedef class obj_type_c;

class object_handle_c;
    object                obj_h;

    virtual function obj_type_c get_obj_type();
        `ZSP_FATAL(("get_obj_type not implemented"));
    endfunction

endclass
