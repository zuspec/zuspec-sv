
class empty_addr_trait_s;

    static function empty_addr_trait_s create_default();
        empty_addr_trait_s ret = new();
        return ret;
    endfunction
endclass
