
class set_c #(type T);
    bit         m_store[T];

    
endclass
