
class pool_c;

endclass